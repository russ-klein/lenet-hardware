module dump;

initial $fsdbDumpvars;

endmodule
